//////////////////////////////////////////////////////////////////////////////////
// Engineer: 		Travis
// 
// Create Date: 	11/13/2020 Wed 16:36
// Filename: 		apb_slv_pkg.svh
// class Name: 		apb_slv_pkg
// Project Name: 	ahb2apb_bridge
// Revision 0.01 - File Created
// Additional Comments:
// -------------------------------------------------------------------------------
//////////////////////////////////////////////////////////////////////////////////
`ifndef APB_SLAVE_ENUM_SV
`define APB_SLAVE_ENUM_SV

    typedef enum {READ, WRITE} kind_t;

`endif
