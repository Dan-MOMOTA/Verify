module queue;
    int j=1,
    q2[$]={3,4},
    q[$]={0,2,5};          //声明队列,并初始化一些元素
    initial begin
        q.insert(1,j);     // 在q队列的第二个元素(排列位置从0开始数)之前插入j,// 队列q变成{0,1,2,5}
        q.insert(3,q2[0]); //在q队列的第四个元素(排列位置从0开始数)之前
        q.insert(4,q2[1]); // 插入队列q2的元素，队列q变成{0,1,2,3,4,5}
        $display(q);
        q.delete(1);       //删除第1个元素(排列位置从0开始数), 队列变成{0,2,3,4,5}
        q.push_front(6);   //在队列前插入6, q队列变成{6,0,2,3,4,5}
        j = q.pop_back;    //把最后一个元素pop出来,赋值给j, j=5, q队列变成{6,0,2,3,4}
        q.push_back(8);    //在队列尾部插入8, q队列变成{6,0,2,3,4,8}
        j = q.pop_front;   //把第一个元素pop出来,赋值给j, j=6, q队列变成{0,2,3,4,8}
        foreach (q[i])
            $display(q[i]);    //打印整个队列
        q.delete();        //删除整个队列
    end
endmodule

//队列的声明使用[$],q[$:其他]：
//把$放在一个范围表达式的左边，那么$代表最小值
//把$放在一个范围表达式的右边，那么$代表最大值