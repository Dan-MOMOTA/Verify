module test_top;

    real a ;
    int  b ;
    real c ;

    initial begin

        a = 14/5;
        b = a;
        c = 14.0/5;

        $display("a = %0f, b = %0d , c = %0f", a, b, c);
    end

endmodule

/*
 *仿真结果
 *a = 2.000000, b = 2, c = 2.800000
 *在Verilog中,实数类型的变量默认是双精度浮点数。当你将一个整数除以另一个整数时,
 *Verilog会执行整数除法,结果将会是一个整数,小数部分会被舍去。因此,14除以5的结果是2,
 *因为它执行的是整数除法。如果你希望得到2.8这个结果,你可以将14或5其中一个转换为实数类型,
 *例如14.0/5或14/5.0。这样除法操作将会执行实数除法，得到正确的结果。
 */
