module test_top;

endmodule
